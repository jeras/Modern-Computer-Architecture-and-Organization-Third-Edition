../../Chapter Files/ALU.vhdl